`timescale 1ns / 1ps

module tb();
	reg clk;
	reg reset;
	
	wire [31:0] WriteData, dataadr;
	wire MemWrite;
	
// instantiate device to be tested
main dut(clk, reset, WriteData, dataadr, MemWrite);

// initialize test
initial
	begin
	reset <= 1; # 22; reset <= 0;
end

// generate clock to sequence tests
always
	begin
	clk <= 1; # 5; 
	clk <= 0; # 5;
end

// check results
always @ (negedge clk)
	begin
		if (MemWrite) begin
		if (dataadr === 84 & WriteData === 7) begin
			$display ("Simulation succeeded");
			$stop;
			
	end else if (dataadr !== 80) begin
				$display ("Simulation failed");
				$stop;
		end
	end
end

endmodule 